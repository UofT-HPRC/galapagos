`timescale 1 ps / 1 ps

module shellTop
   (
    gt_1_ref_clk_n,
    gt_1_ref_clk_p,
    init_clk_n,
    init_clk_p,
    qsfp1_4x_grx_n,
    qsfp1_4x_grx_p,
    qsfp1_4x_gtx_n,
    qsfp1_4x_gtx_p