`timescale 1 ps / 1 ps

module shellTop
   (
    gt_1_ref_clk_n,
    gt_1_ref_clk_p,
    init_clk_n,
    init_clk_p);


  input gt_1_ref_clk_n;
  input gt_1_ref_clk_p;
  input [0:0]init_clk_n;
  input [0:0]init_clk_p;

  wire rstn;
  wire rstn300;
  wire CLK;
  wire CLK300;

  wire gt_1_ref_clk_n;
  wire gt_1_ref_clk_p;
  wire [0:0]init_clk_n;
  wire [0:0]init_clk_p;

